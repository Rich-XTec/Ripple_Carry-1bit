library verilog;
use verilog.vl_types.all;
entity ripple_carry_tb is
end ripple_carry_tb;
